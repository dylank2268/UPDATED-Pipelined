--Dylan Kramer
--5 to 32 decoder

library IEEE;
use IEEE.std_logic_1164.all;
use work.RISCV_types.all;

entity decoder5t32 is
  port (
    DIN  : in  std_logic_vector(4 downto 0);    
    EN: in std_logic;
    Y  : out std_logic_vector(31 downto 0)    
  );
end decoder5t32;

architecture dataflow of decoder5t32 is
begin
	Y <= (others => '0') when EN = '0' else
       "00000000000000000000000000000001" when DIN = "00000" else
       "00000000000000000000000000000010" when DIN = "00001" else
       "00000000000000000000000000000100" when DIN = "00010" else
       "00000000000000000000000000001000" when DIN = "00011" else
       "00000000000000000000000000010000" when DIN = "00100" else
       "00000000000000000000000000100000" when DIN = "00101" else
       "00000000000000000000000001000000" when DIN = "00110" else
       "00000000000000000000000010000000" when DIN = "00111" else
       "00000000000000000000000100000000" when DIN = "01000" else
       "00000000000000000000001000000000" when DIN = "01001" else
       "00000000000000000000010000000000" when DIN = "01010" else
       "00000000000000000000100000000000" when DIN = "01011" else
       "00000000000000000001000000000000" when DIN = "01100" else
       "00000000000000000010000000000000" when DIN = "01101" else
       "00000000000000000100000000000000" when DIN = "01110" else
       "00000000000000001000000000000000" when DIN = "01111" else
       "00000000000000010000000000000000" when DIN = "10000" else
       "00000000000000100000000000000000" when DIN = "10001" else
       "00000000000001000000000000000000" when DIN = "10010" else 
       "00000000000010000000000000000000" when DIN = "10011" else
       "00000000000100000000000000000000" when DIN = "10100" else
       "00000000001000000000000000000000" when DIN = "10101" else
       "00000000010000000000000000000000" when DIN = "10110" else
       "00000000100000000000000000000000" when DIN = "10111" else
       "00000001000000000000000000000000" when DIN = "11000" else
       "00000010000000000000000000000000" when DIN = "11001" else
       "00000100000000000000000000000000" when DIN = "11010" else
       "00001000000000000000000000000000" when DIN = "11011" else
       "00010000000000000000000000000000" when DIN = "11100" else
       "00100000000000000000000000000000" when DIN = "11101" else
       "01000000000000000000000000000000" when DIN = "11110" else
       "10000000000000000000000000000000" when DIN = "11111" else
       (others => '0');  
end dataflow;
